module test_top #(
	parameter INST_MEM_WIDTH = 2
);

